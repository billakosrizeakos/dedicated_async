magic
tech sky130A
magscale 1 2
timestamp 1727860891
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 38824 37584
<< obsm2 >>
rect 938 2139 38530 37573
<< metal3 >>
rect 0 36184 800 36304
rect 0 29656 800 29776
rect 0 23128 800 23248
rect 39200 19864 40000 19984
rect 0 16600 800 16720
rect 0 10072 800 10192
rect 0 3544 800 3664
<< obsm3 >>
rect 798 36384 39200 37569
rect 880 36104 39200 36384
rect 798 29856 39200 36104
rect 880 29576 39200 29856
rect 798 23328 39200 29576
rect 880 23048 39200 23328
rect 798 20064 39200 23048
rect 798 19784 39120 20064
rect 798 16800 39200 19784
rect 880 16520 39200 16800
rect 798 10272 39200 16520
rect 880 9992 39200 10272
rect 798 3744 39200 9992
rect 880 3464 39200 3744
rect 798 2143 39200 3464
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 3544 800 3664 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 39200 19864 40000 19984 6 io_out
port 7 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 8 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 8 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 9 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 472772
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/muller_c_proj/runs/24_10_02_11_20/results/signoff/muller_c_proj.magic.gds
string GDS_START 73796
<< end >>

