magic
tech sky130A
magscale 1 2
timestamp 1728561207
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 38824 37584
<< obsm2 >>
rect 938 2139 38530 37573
<< metal3 >>
rect 0 37000 800 37120
rect 39200 37000 40000 37120
rect 0 36456 800 36576
rect 0 35912 800 36032
rect 0 35368 800 35488
rect 0 34824 800 34944
rect 0 34280 800 34400
rect 0 33736 800 33856
rect 0 33192 800 33312
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 0 31560 800 31680
rect 39200 31288 40000 31408
rect 0 31016 800 31136
rect 0 30472 800 30592
rect 0 29928 800 30048
rect 0 29384 800 29504
rect 0 28840 800 28960
rect 0 28296 800 28416
rect 0 27752 800 27872
rect 0 27208 800 27328
rect 0 26664 800 26784
rect 0 26120 800 26240
rect 0 25576 800 25696
rect 39200 25576 40000 25696
rect 0 25032 800 25152
rect 0 24488 800 24608
rect 0 23944 800 24064
rect 0 23400 800 23520
rect 0 22856 800 22976
rect 0 22312 800 22432
rect 0 21768 800 21888
rect 0 21224 800 21344
rect 0 20680 800 20800
rect 0 20136 800 20256
rect 39200 19864 40000 19984
rect 0 19592 800 19712
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 39200 14152 40000 14272
rect 0 13608 800 13728
rect 0 13064 800 13184
rect 0 12520 800 12640
rect 0 11976 800 12096
rect 0 11432 800 11552
rect 0 10888 800 11008
rect 0 10344 800 10464
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8712 800 8832
rect 39200 8440 40000 8560
rect 0 8168 800 8288
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 0 6536 800 6656
rect 0 5992 800 6112
rect 0 5448 800 5568
rect 0 4904 800 5024
rect 0 4360 800 4480
rect 0 3816 800 3936
rect 0 3272 800 3392
rect 0 2728 800 2848
rect 39200 2728 40000 2848
<< obsm3 >>
rect 798 37200 39200 37569
rect 880 36920 39120 37200
rect 798 36656 39200 36920
rect 880 36376 39200 36656
rect 798 36112 39200 36376
rect 880 35832 39200 36112
rect 798 35568 39200 35832
rect 880 35288 39200 35568
rect 798 35024 39200 35288
rect 880 34744 39200 35024
rect 798 34480 39200 34744
rect 880 34200 39200 34480
rect 798 33936 39200 34200
rect 880 33656 39200 33936
rect 798 33392 39200 33656
rect 880 33112 39200 33392
rect 798 32848 39200 33112
rect 880 32568 39200 32848
rect 798 32304 39200 32568
rect 880 32024 39200 32304
rect 798 31760 39200 32024
rect 880 31488 39200 31760
rect 880 31480 39120 31488
rect 798 31216 39120 31480
rect 880 31208 39120 31216
rect 880 30936 39200 31208
rect 798 30672 39200 30936
rect 880 30392 39200 30672
rect 798 30128 39200 30392
rect 880 29848 39200 30128
rect 798 29584 39200 29848
rect 880 29304 39200 29584
rect 798 29040 39200 29304
rect 880 28760 39200 29040
rect 798 28496 39200 28760
rect 880 28216 39200 28496
rect 798 27952 39200 28216
rect 880 27672 39200 27952
rect 798 27408 39200 27672
rect 880 27128 39200 27408
rect 798 26864 39200 27128
rect 880 26584 39200 26864
rect 798 26320 39200 26584
rect 880 26040 39200 26320
rect 798 25776 39200 26040
rect 880 25496 39120 25776
rect 798 25232 39200 25496
rect 880 24952 39200 25232
rect 798 24688 39200 24952
rect 880 24408 39200 24688
rect 798 24144 39200 24408
rect 880 23864 39200 24144
rect 798 23600 39200 23864
rect 880 23320 39200 23600
rect 798 23056 39200 23320
rect 880 22776 39200 23056
rect 798 22512 39200 22776
rect 880 22232 39200 22512
rect 798 21968 39200 22232
rect 880 21688 39200 21968
rect 798 21424 39200 21688
rect 880 21144 39200 21424
rect 798 20880 39200 21144
rect 880 20600 39200 20880
rect 798 20336 39200 20600
rect 880 20064 39200 20336
rect 880 20056 39120 20064
rect 798 19792 39120 20056
rect 880 19784 39120 19792
rect 880 19512 39200 19784
rect 798 19248 39200 19512
rect 880 18968 39200 19248
rect 798 18704 39200 18968
rect 880 18424 39200 18704
rect 798 18160 39200 18424
rect 880 17880 39200 18160
rect 798 17616 39200 17880
rect 880 17336 39200 17616
rect 798 17072 39200 17336
rect 880 16792 39200 17072
rect 798 16528 39200 16792
rect 880 16248 39200 16528
rect 798 15984 39200 16248
rect 880 15704 39200 15984
rect 798 15440 39200 15704
rect 880 15160 39200 15440
rect 798 14896 39200 15160
rect 880 14616 39200 14896
rect 798 14352 39200 14616
rect 880 14072 39120 14352
rect 798 13808 39200 14072
rect 880 13528 39200 13808
rect 798 13264 39200 13528
rect 880 12984 39200 13264
rect 798 12720 39200 12984
rect 880 12440 39200 12720
rect 798 12176 39200 12440
rect 880 11896 39200 12176
rect 798 11632 39200 11896
rect 880 11352 39200 11632
rect 798 11088 39200 11352
rect 880 10808 39200 11088
rect 798 10544 39200 10808
rect 880 10264 39200 10544
rect 798 10000 39200 10264
rect 880 9720 39200 10000
rect 798 9456 39200 9720
rect 880 9176 39200 9456
rect 798 8912 39200 9176
rect 880 8640 39200 8912
rect 880 8632 39120 8640
rect 798 8368 39120 8632
rect 880 8360 39120 8368
rect 880 8088 39200 8360
rect 798 7824 39200 8088
rect 880 7544 39200 7824
rect 798 7280 39200 7544
rect 880 7000 39200 7280
rect 798 6736 39200 7000
rect 880 6456 39200 6736
rect 798 6192 39200 6456
rect 880 5912 39200 6192
rect 798 5648 39200 5912
rect 880 5368 39200 5648
rect 798 5104 39200 5368
rect 880 4824 39200 5104
rect 798 4560 39200 4824
rect 880 4280 39200 4560
rect 798 4016 39200 4280
rect 880 3736 39200 4016
rect 798 3472 39200 3736
rect 880 3192 39200 3472
rect 798 2928 39200 3192
rect 880 2648 39120 2928
rect 798 2143 39200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 2728 800 2848 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 io_in[38]
port 32 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 io_in[39]
port 33 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 io_in[3]
port 34 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[40]
port 35 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 io_in[41]
port 36 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 io_in[42]
port 37 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 io_in[43]
port 38 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 io_in[44]
port 39 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_in[45]
port 40 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 io_in[46]
port 41 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 io_in[47]
port 42 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[48]
port 43 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 io_in[49]
port 44 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 io_in[4]
port 45 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_in[50]
port 46 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 io_in[51]
port 47 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 io_in[52]
port 48 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 io_in[53]
port 49 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 io_in[54]
port 50 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 io_in[55]
port 51 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 io_in[56]
port 52 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 io_in[57]
port 53 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 io_in[58]
port 54 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 io_in[59]
port 55 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_in[5]
port 56 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_in[60]
port 57 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 io_in[61]
port 58 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 io_in[62]
port 59 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 io_in[63]
port 60 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 io_in[6]
port 61 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 io_in[7]
port 62 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 io_in[8]
port 63 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 io_in[9]
port 64 nsew signal input
rlabel metal3 s 39200 2728 40000 2848 6 io_out[0]
port 65 nsew signal output
rlabel metal3 s 39200 8440 40000 8560 6 io_out[1]
port 66 nsew signal output
rlabel metal3 s 39200 14152 40000 14272 6 io_out[2]
port 67 nsew signal output
rlabel metal3 s 39200 19864 40000 19984 6 io_out[3]
port 68 nsew signal output
rlabel metal3 s 39200 25576 40000 25696 6 io_out[4]
port 69 nsew signal output
rlabel metal3 s 39200 31288 40000 31408 6 io_out[5]
port 70 nsew signal output
rlabel metal3 s 39200 37000 40000 37120 6 valid
port 71 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 72 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 72 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 73 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 877744
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/encoder_proj/runs/24_10_10_13_52/results/signoff/encoder_proj.magic.gds
string GDS_START 164798
<< end >>

