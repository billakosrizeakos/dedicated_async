VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder_proj
  CLASS BLOCK ;
  FOREIGN decoder_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END enable
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_in[5]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 200.000 14.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.840 200.000 41.440 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 43.560 200.000 44.160 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.280 200.000 46.880 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.000 200.000 49.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.720 200.000 52.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 200.000 55.040 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 57.160 200.000 57.760 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 59.880 200.000 60.480 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 62.600 200.000 63.200 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 65.320 200.000 65.920 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 16.360 200.000 16.960 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.040 200.000 68.640 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.760 200.000 71.360 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 73.480 200.000 74.080 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 76.200 200.000 76.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.920 200.000 79.520 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 84.360 200.000 84.960 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.080 200.000 87.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.800 200.000 90.400 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 92.520 200.000 93.120 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 19.080 200.000 19.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 97.960 200.000 98.560 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 100.680 200.000 101.280 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 103.400 200.000 104.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 106.120 200.000 106.720 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 200.000 109.440 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 111.560 200.000 112.160 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.280 200.000 114.880 ;
    END
  END io_out[37]
  PIN io_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 117.000 200.000 117.600 ;
    END
  END io_out[38]
  PIN io_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.720 200.000 120.320 ;
    END
  END io_out[39]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 21.800 200.000 22.400 ;
    END
  END io_out[3]
  PIN io_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 122.440 200.000 123.040 ;
    END
  END io_out[40]
  PIN io_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.160 200.000 125.760 ;
    END
  END io_out[41]
  PIN io_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 200.000 128.480 ;
    END
  END io_out[42]
  PIN io_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 130.600 200.000 131.200 ;
    END
  END io_out[43]
  PIN io_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 133.320 200.000 133.920 ;
    END
  END io_out[44]
  PIN io_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 200.000 136.640 ;
    END
  END io_out[45]
  PIN io_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 138.760 200.000 139.360 ;
    END
  END io_out[46]
  PIN io_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 200.000 142.080 ;
    END
  END io_out[47]
  PIN io_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 144.200 200.000 144.800 ;
    END
  END io_out[48]
  PIN io_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 146.920 200.000 147.520 ;
    END
  END io_out[49]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 24.520 200.000 25.120 ;
    END
  END io_out[4]
  PIN io_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 149.640 200.000 150.240 ;
    END
  END io_out[50]
  PIN io_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END io_out[51]
  PIN io_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 200.000 155.680 ;
    END
  END io_out[52]
  PIN io_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.800 200.000 158.400 ;
    END
  END io_out[53]
  PIN io_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 160.520 200.000 161.120 ;
    END
  END io_out[54]
  PIN io_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END io_out[55]
  PIN io_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 200.000 166.560 ;
    END
  END io_out[56]
  PIN io_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END io_out[57]
  PIN io_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 171.400 200.000 172.000 ;
    END
  END io_out[58]
  PIN io_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.120 200.000 174.720 ;
    END
  END io_out[59]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.240 200.000 27.840 ;
    END
  END io_out[5]
  PIN io_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END io_out[60]
  PIN io_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 200.000 180.160 ;
    END
  END io_out[61]
  PIN io_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 182.280 200.000 182.880 ;
    END
  END io_out[62]
  PIN io_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.000 200.000 185.600 ;
    END
  END io_out[63]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.960 200.000 30.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.680 200.000 33.280 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 35.400 200.000 36.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 38.120 200.000 38.720 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 199.570 187.920 ;
      LAYER met2 ;
        RECT 4.690 10.695 199.540 187.865 ;
      LAYER met3 ;
        RECT 3.990 186.000 196.000 187.845 ;
        RECT 4.400 184.600 195.600 186.000 ;
        RECT 3.990 183.280 196.000 184.600 ;
        RECT 3.990 181.880 195.600 183.280 ;
        RECT 3.990 180.560 196.000 181.880 ;
        RECT 3.990 179.160 195.600 180.560 ;
        RECT 3.990 177.840 196.000 179.160 ;
        RECT 3.990 176.440 195.600 177.840 ;
        RECT 3.990 175.120 196.000 176.440 ;
        RECT 3.990 173.720 195.600 175.120 ;
        RECT 3.990 172.400 196.000 173.720 ;
        RECT 3.990 171.000 195.600 172.400 ;
        RECT 3.990 169.680 196.000 171.000 ;
        RECT 3.990 168.280 195.600 169.680 ;
        RECT 3.990 166.960 196.000 168.280 ;
        RECT 3.990 165.560 195.600 166.960 ;
        RECT 3.990 164.240 196.000 165.560 ;
        RECT 3.990 162.840 195.600 164.240 ;
        RECT 3.990 161.520 196.000 162.840 ;
        RECT 3.990 160.120 195.600 161.520 ;
        RECT 3.990 158.800 196.000 160.120 ;
        RECT 3.990 157.440 195.600 158.800 ;
        RECT 4.400 157.400 195.600 157.440 ;
        RECT 4.400 156.080 196.000 157.400 ;
        RECT 4.400 156.040 195.600 156.080 ;
        RECT 3.990 154.680 195.600 156.040 ;
        RECT 3.990 153.360 196.000 154.680 ;
        RECT 3.990 151.960 195.600 153.360 ;
        RECT 3.990 150.640 196.000 151.960 ;
        RECT 3.990 149.240 195.600 150.640 ;
        RECT 3.990 147.920 196.000 149.240 ;
        RECT 3.990 146.520 195.600 147.920 ;
        RECT 3.990 145.200 196.000 146.520 ;
        RECT 3.990 143.800 195.600 145.200 ;
        RECT 3.990 142.480 196.000 143.800 ;
        RECT 3.990 141.080 195.600 142.480 ;
        RECT 3.990 139.760 196.000 141.080 ;
        RECT 3.990 138.360 195.600 139.760 ;
        RECT 3.990 137.040 196.000 138.360 ;
        RECT 3.990 135.640 195.600 137.040 ;
        RECT 3.990 134.320 196.000 135.640 ;
        RECT 3.990 132.920 195.600 134.320 ;
        RECT 3.990 131.600 196.000 132.920 ;
        RECT 3.990 130.200 195.600 131.600 ;
        RECT 3.990 128.880 196.000 130.200 ;
        RECT 4.400 127.480 195.600 128.880 ;
        RECT 3.990 126.160 196.000 127.480 ;
        RECT 3.990 124.760 195.600 126.160 ;
        RECT 3.990 123.440 196.000 124.760 ;
        RECT 3.990 122.040 195.600 123.440 ;
        RECT 3.990 120.720 196.000 122.040 ;
        RECT 3.990 119.320 195.600 120.720 ;
        RECT 3.990 118.000 196.000 119.320 ;
        RECT 3.990 116.600 195.600 118.000 ;
        RECT 3.990 115.280 196.000 116.600 ;
        RECT 3.990 113.880 195.600 115.280 ;
        RECT 3.990 112.560 196.000 113.880 ;
        RECT 3.990 111.160 195.600 112.560 ;
        RECT 3.990 109.840 196.000 111.160 ;
        RECT 3.990 108.440 195.600 109.840 ;
        RECT 3.990 107.120 196.000 108.440 ;
        RECT 3.990 105.720 195.600 107.120 ;
        RECT 3.990 104.400 196.000 105.720 ;
        RECT 3.990 103.000 195.600 104.400 ;
        RECT 3.990 101.680 196.000 103.000 ;
        RECT 3.990 100.320 195.600 101.680 ;
        RECT 4.400 100.280 195.600 100.320 ;
        RECT 4.400 98.960 196.000 100.280 ;
        RECT 4.400 98.920 195.600 98.960 ;
        RECT 3.990 97.560 195.600 98.920 ;
        RECT 3.990 96.240 196.000 97.560 ;
        RECT 3.990 94.840 195.600 96.240 ;
        RECT 3.990 93.520 196.000 94.840 ;
        RECT 3.990 92.120 195.600 93.520 ;
        RECT 3.990 90.800 196.000 92.120 ;
        RECT 3.990 89.400 195.600 90.800 ;
        RECT 3.990 88.080 196.000 89.400 ;
        RECT 3.990 86.680 195.600 88.080 ;
        RECT 3.990 85.360 196.000 86.680 ;
        RECT 3.990 83.960 195.600 85.360 ;
        RECT 3.990 82.640 196.000 83.960 ;
        RECT 3.990 81.240 195.600 82.640 ;
        RECT 3.990 79.920 196.000 81.240 ;
        RECT 3.990 78.520 195.600 79.920 ;
        RECT 3.990 77.200 196.000 78.520 ;
        RECT 3.990 75.800 195.600 77.200 ;
        RECT 3.990 74.480 196.000 75.800 ;
        RECT 3.990 73.080 195.600 74.480 ;
        RECT 3.990 71.760 196.000 73.080 ;
        RECT 4.400 70.360 195.600 71.760 ;
        RECT 3.990 69.040 196.000 70.360 ;
        RECT 3.990 67.640 195.600 69.040 ;
        RECT 3.990 66.320 196.000 67.640 ;
        RECT 3.990 64.920 195.600 66.320 ;
        RECT 3.990 63.600 196.000 64.920 ;
        RECT 3.990 62.200 195.600 63.600 ;
        RECT 3.990 60.880 196.000 62.200 ;
        RECT 3.990 59.480 195.600 60.880 ;
        RECT 3.990 58.160 196.000 59.480 ;
        RECT 3.990 56.760 195.600 58.160 ;
        RECT 3.990 55.440 196.000 56.760 ;
        RECT 3.990 54.040 195.600 55.440 ;
        RECT 3.990 52.720 196.000 54.040 ;
        RECT 3.990 51.320 195.600 52.720 ;
        RECT 3.990 50.000 196.000 51.320 ;
        RECT 3.990 48.600 195.600 50.000 ;
        RECT 3.990 47.280 196.000 48.600 ;
        RECT 3.990 45.880 195.600 47.280 ;
        RECT 3.990 44.560 196.000 45.880 ;
        RECT 3.990 43.200 195.600 44.560 ;
        RECT 4.400 43.160 195.600 43.200 ;
        RECT 4.400 41.840 196.000 43.160 ;
        RECT 4.400 41.800 195.600 41.840 ;
        RECT 3.990 40.440 195.600 41.800 ;
        RECT 3.990 39.120 196.000 40.440 ;
        RECT 3.990 37.720 195.600 39.120 ;
        RECT 3.990 36.400 196.000 37.720 ;
        RECT 3.990 35.000 195.600 36.400 ;
        RECT 3.990 33.680 196.000 35.000 ;
        RECT 3.990 32.280 195.600 33.680 ;
        RECT 3.990 30.960 196.000 32.280 ;
        RECT 3.990 29.560 195.600 30.960 ;
        RECT 3.990 28.240 196.000 29.560 ;
        RECT 3.990 26.840 195.600 28.240 ;
        RECT 3.990 25.520 196.000 26.840 ;
        RECT 3.990 24.120 195.600 25.520 ;
        RECT 3.990 22.800 196.000 24.120 ;
        RECT 3.990 21.400 195.600 22.800 ;
        RECT 3.990 20.080 196.000 21.400 ;
        RECT 3.990 18.680 195.600 20.080 ;
        RECT 3.990 17.360 196.000 18.680 ;
        RECT 3.990 15.960 195.600 17.360 ;
        RECT 3.990 14.640 196.000 15.960 ;
        RECT 4.400 13.240 195.600 14.640 ;
        RECT 3.990 10.715 196.000 13.240 ;
  END
END decoder_proj
END LIBRARY

