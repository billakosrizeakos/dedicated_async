magic
tech sky130A
magscale 1 2
timestamp 1728465731
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 38824 37584
<< obsm2 >>
rect 938 2139 38530 37573
<< metal3 >>
rect 0 33192 800 33312
rect 39200 33192 40000 33312
rect 0 19864 800 19984
rect 39200 19864 40000 19984
rect 0 6536 800 6656
rect 39200 6536 40000 6656
<< obsm3 >>
rect 800 33392 39200 37569
rect 880 33112 39120 33392
rect 800 20064 39200 33112
rect 880 19784 39120 20064
rect 800 6736 39200 19784
rect 880 6456 39120 6736
rect 800 2143 39200 6456
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 6536 800 6656 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 39200 6536 40000 6656 6 io_out[0]
port 4 nsew signal output
rlabel metal3 s 39200 19864 40000 19984 6 io_out[1]
port 5 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 io_out[2]
port 6 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 473328
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/arbiter_proj/runs/24_10_09_11_21/results/signoff/arbiter_proj.magic.gds
string GDS_START 59116
<< end >>

