VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO arbiter_cell_two_bits_fc
  CLASS BLOCK ;
  FOREIGN arbiter_cell_two_bits_fc ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END GND
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END VDD
  PIN g0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END g0
  PIN g1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END g1
  PIN gc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 200.000 148.880 ;
    END
  END gc
  PIN r0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END r0
  PIN r1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END r1
  PIN rc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.000 200.000 49.600 ;
    END
  END rc
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.510 187.920 ;
      LAYER met2 ;
        RECT 4.690 10.695 194.490 187.865 ;
      LAYER met3 ;
        RECT 3.990 173.760 196.000 187.845 ;
        RECT 4.400 172.360 196.000 173.760 ;
        RECT 3.990 149.280 196.000 172.360 ;
        RECT 3.990 147.880 195.600 149.280 ;
        RECT 3.990 124.800 196.000 147.880 ;
        RECT 4.400 123.400 196.000 124.800 ;
        RECT 3.990 75.840 196.000 123.400 ;
        RECT 4.400 74.440 196.000 75.840 ;
        RECT 3.990 50.000 196.000 74.440 ;
        RECT 3.990 48.600 195.600 50.000 ;
        RECT 3.990 26.880 196.000 48.600 ;
        RECT 4.400 25.480 196.000 26.880 ;
        RECT 3.990 10.715 196.000 25.480 ;
  END
END arbiter_cell_two_bits_fc
END LIBRARY

