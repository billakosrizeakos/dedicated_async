magic
tech sky130A
magscale 1 2
timestamp 1727860641
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 39914 37584
<< obsm2 >>
rect 938 2139 39908 37573
<< metal3 >>
rect 0 37000 800 37120
rect 39200 37000 40000 37120
rect 39200 36456 40000 36576
rect 39200 35912 40000 36032
rect 39200 35368 40000 35488
rect 39200 34824 40000 34944
rect 39200 34280 40000 34400
rect 39200 33736 40000 33856
rect 39200 33192 40000 33312
rect 39200 32648 40000 32768
rect 39200 32104 40000 32224
rect 39200 31560 40000 31680
rect 0 31288 800 31408
rect 39200 31016 40000 31136
rect 39200 30472 40000 30592
rect 39200 29928 40000 30048
rect 39200 29384 40000 29504
rect 39200 28840 40000 28960
rect 39200 28296 40000 28416
rect 39200 27752 40000 27872
rect 39200 27208 40000 27328
rect 39200 26664 40000 26784
rect 39200 26120 40000 26240
rect 0 25576 800 25696
rect 39200 25576 40000 25696
rect 39200 25032 40000 25152
rect 39200 24488 40000 24608
rect 39200 23944 40000 24064
rect 39200 23400 40000 23520
rect 39200 22856 40000 22976
rect 39200 22312 40000 22432
rect 39200 21768 40000 21888
rect 39200 21224 40000 21344
rect 39200 20680 40000 20800
rect 39200 20136 40000 20256
rect 0 19864 800 19984
rect 39200 19592 40000 19712
rect 39200 19048 40000 19168
rect 39200 18504 40000 18624
rect 39200 17960 40000 18080
rect 39200 17416 40000 17536
rect 39200 16872 40000 16992
rect 39200 16328 40000 16448
rect 39200 15784 40000 15904
rect 39200 15240 40000 15360
rect 39200 14696 40000 14816
rect 0 14152 800 14272
rect 39200 14152 40000 14272
rect 39200 13608 40000 13728
rect 39200 13064 40000 13184
rect 39200 12520 40000 12640
rect 39200 11976 40000 12096
rect 39200 11432 40000 11552
rect 39200 10888 40000 11008
rect 39200 10344 40000 10464
rect 39200 9800 40000 9920
rect 39200 9256 40000 9376
rect 39200 8712 40000 8832
rect 0 8440 800 8560
rect 39200 8168 40000 8288
rect 39200 7624 40000 7744
rect 39200 7080 40000 7200
rect 39200 6536 40000 6656
rect 39200 5992 40000 6112
rect 39200 5448 40000 5568
rect 39200 4904 40000 5024
rect 39200 4360 40000 4480
rect 39200 3816 40000 3936
rect 39200 3272 40000 3392
rect 0 2728 800 2848
rect 39200 2728 40000 2848
<< obsm3 >>
rect 798 37200 39200 37569
rect 880 36920 39120 37200
rect 798 36656 39200 36920
rect 798 36376 39120 36656
rect 798 36112 39200 36376
rect 798 35832 39120 36112
rect 798 35568 39200 35832
rect 798 35288 39120 35568
rect 798 35024 39200 35288
rect 798 34744 39120 35024
rect 798 34480 39200 34744
rect 798 34200 39120 34480
rect 798 33936 39200 34200
rect 798 33656 39120 33936
rect 798 33392 39200 33656
rect 798 33112 39120 33392
rect 798 32848 39200 33112
rect 798 32568 39120 32848
rect 798 32304 39200 32568
rect 798 32024 39120 32304
rect 798 31760 39200 32024
rect 798 31488 39120 31760
rect 880 31480 39120 31488
rect 880 31216 39200 31480
rect 880 31208 39120 31216
rect 798 30936 39120 31208
rect 798 30672 39200 30936
rect 798 30392 39120 30672
rect 798 30128 39200 30392
rect 798 29848 39120 30128
rect 798 29584 39200 29848
rect 798 29304 39120 29584
rect 798 29040 39200 29304
rect 798 28760 39120 29040
rect 798 28496 39200 28760
rect 798 28216 39120 28496
rect 798 27952 39200 28216
rect 798 27672 39120 27952
rect 798 27408 39200 27672
rect 798 27128 39120 27408
rect 798 26864 39200 27128
rect 798 26584 39120 26864
rect 798 26320 39200 26584
rect 798 26040 39120 26320
rect 798 25776 39200 26040
rect 880 25496 39120 25776
rect 798 25232 39200 25496
rect 798 24952 39120 25232
rect 798 24688 39200 24952
rect 798 24408 39120 24688
rect 798 24144 39200 24408
rect 798 23864 39120 24144
rect 798 23600 39200 23864
rect 798 23320 39120 23600
rect 798 23056 39200 23320
rect 798 22776 39120 23056
rect 798 22512 39200 22776
rect 798 22232 39120 22512
rect 798 21968 39200 22232
rect 798 21688 39120 21968
rect 798 21424 39200 21688
rect 798 21144 39120 21424
rect 798 20880 39200 21144
rect 798 20600 39120 20880
rect 798 20336 39200 20600
rect 798 20064 39120 20336
rect 880 20056 39120 20064
rect 880 19792 39200 20056
rect 880 19784 39120 19792
rect 798 19512 39120 19784
rect 798 19248 39200 19512
rect 798 18968 39120 19248
rect 798 18704 39200 18968
rect 798 18424 39120 18704
rect 798 18160 39200 18424
rect 798 17880 39120 18160
rect 798 17616 39200 17880
rect 798 17336 39120 17616
rect 798 17072 39200 17336
rect 798 16792 39120 17072
rect 798 16528 39200 16792
rect 798 16248 39120 16528
rect 798 15984 39200 16248
rect 798 15704 39120 15984
rect 798 15440 39200 15704
rect 798 15160 39120 15440
rect 798 14896 39200 15160
rect 798 14616 39120 14896
rect 798 14352 39200 14616
rect 880 14072 39120 14352
rect 798 13808 39200 14072
rect 798 13528 39120 13808
rect 798 13264 39200 13528
rect 798 12984 39120 13264
rect 798 12720 39200 12984
rect 798 12440 39120 12720
rect 798 12176 39200 12440
rect 798 11896 39120 12176
rect 798 11632 39200 11896
rect 798 11352 39120 11632
rect 798 11088 39200 11352
rect 798 10808 39120 11088
rect 798 10544 39200 10808
rect 798 10264 39120 10544
rect 798 10000 39200 10264
rect 798 9720 39120 10000
rect 798 9456 39200 9720
rect 798 9176 39120 9456
rect 798 8912 39200 9176
rect 798 8640 39120 8912
rect 880 8632 39120 8640
rect 880 8368 39200 8632
rect 880 8360 39120 8368
rect 798 8088 39120 8360
rect 798 7824 39200 8088
rect 798 7544 39120 7824
rect 798 7280 39200 7544
rect 798 7000 39120 7280
rect 798 6736 39200 7000
rect 798 6456 39120 6736
rect 798 6192 39200 6456
rect 798 5912 39120 6192
rect 798 5648 39200 5912
rect 798 5368 39120 5648
rect 798 5104 39200 5368
rect 798 4824 39120 5104
rect 798 4560 39200 4824
rect 798 4280 39120 4560
rect 798 4016 39200 4280
rect 798 3736 39120 4016
rect 798 3472 39200 3736
rect 798 3192 39120 3472
rect 798 2928 39200 3192
rect 880 2648 39120 2928
rect 798 2143 39200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 37000 800 37120 6 enable
port 1 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 39200 2728 40000 2848 6 io_out[0]
port 8 nsew signal output
rlabel metal3 s 39200 8168 40000 8288 6 io_out[10]
port 9 nsew signal output
rlabel metal3 s 39200 8712 40000 8832 6 io_out[11]
port 10 nsew signal output
rlabel metal3 s 39200 9256 40000 9376 6 io_out[12]
port 11 nsew signal output
rlabel metal3 s 39200 9800 40000 9920 6 io_out[13]
port 12 nsew signal output
rlabel metal3 s 39200 10344 40000 10464 6 io_out[14]
port 13 nsew signal output
rlabel metal3 s 39200 10888 40000 11008 6 io_out[15]
port 14 nsew signal output
rlabel metal3 s 39200 11432 40000 11552 6 io_out[16]
port 15 nsew signal output
rlabel metal3 s 39200 11976 40000 12096 6 io_out[17]
port 16 nsew signal output
rlabel metal3 s 39200 12520 40000 12640 6 io_out[18]
port 17 nsew signal output
rlabel metal3 s 39200 13064 40000 13184 6 io_out[19]
port 18 nsew signal output
rlabel metal3 s 39200 3272 40000 3392 6 io_out[1]
port 19 nsew signal output
rlabel metal3 s 39200 13608 40000 13728 6 io_out[20]
port 20 nsew signal output
rlabel metal3 s 39200 14152 40000 14272 6 io_out[21]
port 21 nsew signal output
rlabel metal3 s 39200 14696 40000 14816 6 io_out[22]
port 22 nsew signal output
rlabel metal3 s 39200 15240 40000 15360 6 io_out[23]
port 23 nsew signal output
rlabel metal3 s 39200 15784 40000 15904 6 io_out[24]
port 24 nsew signal output
rlabel metal3 s 39200 16328 40000 16448 6 io_out[25]
port 25 nsew signal output
rlabel metal3 s 39200 16872 40000 16992 6 io_out[26]
port 26 nsew signal output
rlabel metal3 s 39200 17416 40000 17536 6 io_out[27]
port 27 nsew signal output
rlabel metal3 s 39200 17960 40000 18080 6 io_out[28]
port 28 nsew signal output
rlabel metal3 s 39200 18504 40000 18624 6 io_out[29]
port 29 nsew signal output
rlabel metal3 s 39200 3816 40000 3936 6 io_out[2]
port 30 nsew signal output
rlabel metal3 s 39200 19048 40000 19168 6 io_out[30]
port 31 nsew signal output
rlabel metal3 s 39200 19592 40000 19712 6 io_out[31]
port 32 nsew signal output
rlabel metal3 s 39200 20136 40000 20256 6 io_out[32]
port 33 nsew signal output
rlabel metal3 s 39200 20680 40000 20800 6 io_out[33]
port 34 nsew signal output
rlabel metal3 s 39200 21224 40000 21344 6 io_out[34]
port 35 nsew signal output
rlabel metal3 s 39200 21768 40000 21888 6 io_out[35]
port 36 nsew signal output
rlabel metal3 s 39200 22312 40000 22432 6 io_out[36]
port 37 nsew signal output
rlabel metal3 s 39200 22856 40000 22976 6 io_out[37]
port 38 nsew signal output
rlabel metal3 s 39200 23400 40000 23520 6 io_out[38]
port 39 nsew signal output
rlabel metal3 s 39200 23944 40000 24064 6 io_out[39]
port 40 nsew signal output
rlabel metal3 s 39200 4360 40000 4480 6 io_out[3]
port 41 nsew signal output
rlabel metal3 s 39200 24488 40000 24608 6 io_out[40]
port 42 nsew signal output
rlabel metal3 s 39200 25032 40000 25152 6 io_out[41]
port 43 nsew signal output
rlabel metal3 s 39200 25576 40000 25696 6 io_out[42]
port 44 nsew signal output
rlabel metal3 s 39200 26120 40000 26240 6 io_out[43]
port 45 nsew signal output
rlabel metal3 s 39200 26664 40000 26784 6 io_out[44]
port 46 nsew signal output
rlabel metal3 s 39200 27208 40000 27328 6 io_out[45]
port 47 nsew signal output
rlabel metal3 s 39200 27752 40000 27872 6 io_out[46]
port 48 nsew signal output
rlabel metal3 s 39200 28296 40000 28416 6 io_out[47]
port 49 nsew signal output
rlabel metal3 s 39200 28840 40000 28960 6 io_out[48]
port 50 nsew signal output
rlabel metal3 s 39200 29384 40000 29504 6 io_out[49]
port 51 nsew signal output
rlabel metal3 s 39200 4904 40000 5024 6 io_out[4]
port 52 nsew signal output
rlabel metal3 s 39200 29928 40000 30048 6 io_out[50]
port 53 nsew signal output
rlabel metal3 s 39200 30472 40000 30592 6 io_out[51]
port 54 nsew signal output
rlabel metal3 s 39200 31016 40000 31136 6 io_out[52]
port 55 nsew signal output
rlabel metal3 s 39200 31560 40000 31680 6 io_out[53]
port 56 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 io_out[54]
port 57 nsew signal output
rlabel metal3 s 39200 32648 40000 32768 6 io_out[55]
port 58 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 io_out[56]
port 59 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 io_out[57]
port 60 nsew signal output
rlabel metal3 s 39200 34280 40000 34400 6 io_out[58]
port 61 nsew signal output
rlabel metal3 s 39200 34824 40000 34944 6 io_out[59]
port 62 nsew signal output
rlabel metal3 s 39200 5448 40000 5568 6 io_out[5]
port 63 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 io_out[60]
port 64 nsew signal output
rlabel metal3 s 39200 35912 40000 36032 6 io_out[61]
port 65 nsew signal output
rlabel metal3 s 39200 36456 40000 36576 6 io_out[62]
port 66 nsew signal output
rlabel metal3 s 39200 37000 40000 37120 6 io_out[63]
port 67 nsew signal output
rlabel metal3 s 39200 5992 40000 6112 6 io_out[6]
port 68 nsew signal output
rlabel metal3 s 39200 6536 40000 6656 6 io_out[7]
port 69 nsew signal output
rlabel metal3 s 39200 7080 40000 7200 6 io_out[8]
port 70 nsew signal output
rlabel metal3 s 39200 7624 40000 7744 6 io_out[9]
port 71 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 72 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 72 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 73 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 887852
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/decoder_proj/runs/24_10_02_11_16/results/signoff/decoder_proj.magic.gds
string GDS_START 148808
<< end >>

