* NGSPICE file created from arbiter_cell_two_bits_fc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt arbiter_cell_two_bits_fc GND VDD g0 g1 gc r0 r1 rc GND_uq0 VDD_uq0
XTAP_188 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_49_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_27_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XANTENNA_x2_B x6/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_38_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_507 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_529 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_518 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_12_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_348 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_189 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_63_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx1 x7/Y x6/X GND GND VDD VDD x8/D sky130_fd_sc_hd__nand2_1
XFILLER_0_19_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_59_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XTAP_519 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_35_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_18 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_38_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_349 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_305 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_179 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_23_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xx2 x2/A x6/A GND GND VDD VDD x7/A sky130_fd_sc_hd__or2_1
XFILLER_0_63_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_19_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_509 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_339 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_169 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_46_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xx3 x4/X x9/A GND GND VDD VDD x3/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_20 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_34_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_307 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_58_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_137 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_159 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_490 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx4 x7/Y x7/Y x7/Y x7/Y GND GND VDD VDD x4/X sky130_fd_sc_hd__or4_1
XFILLER_0_39_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_42_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_21_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_308 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_25_3 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_35_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_138 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_54 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_57_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_17_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_491 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx5 x6/A GND GND VDD VDD x9/A sky130_fd_sc_hd__inv_1
XFILLER_0_54_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_33_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_309 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_120 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_139 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_22 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_32_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_492 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx6 x6/A x6/B GND GND VDD VDD x6/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_61_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_121 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_110 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_34 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_25_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_493 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xx7 x7/A x8/D GND GND VDD VDD x7/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_290 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_100 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_122 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_111 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_40_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_494 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx8 x8/D x8/D x8/D x8/D GND GND VDD VDD x9/B sky130_fd_sc_hd__or4_1
XFILLER_0_54_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_280 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_34_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_123 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_112 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_101 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_14 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_27_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_40_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_495 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx9 x9/A x9/B GND GND VDD VDD x9/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_270 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_124 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_113 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_102 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_441 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_496 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_260 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_125 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_114 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_103 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_63_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_475 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_497 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_250 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_35_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_25_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_397 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_7_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_30_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_126 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_115 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_104 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_34_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_389 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_63_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_498 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_240 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xinput1 gc GND GND VDD VDD x6/A sky130_fd_sc_hd__buf_2
XFILLER_0_46_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XANTENNA_x5_A x6/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_116 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_105 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_127 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_27_18 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_57_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_31_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_400 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_499 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_230 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_252 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_9_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_60_9 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xinput2 r0 GND GND VDD VDD x2/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_128 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_117 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_106 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_31_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_423 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_489 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_220 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_286 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_18_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xinput3 r1 GND GND VDD VDD x6/B sky130_fd_sc_hd__buf_1
XFILLER_0_61_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_57_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_43_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_129 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_118 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_107 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_457 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_479 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XTAP_210 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_29_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_55_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_50_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_20 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_32_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_61_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_119 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_108 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_469 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XTAP_200 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_32 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_48_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_35_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_459 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_201 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_44 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_90 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_56_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_405 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_449 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_202 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XTAP_268 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_91 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_80 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_6 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_439 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_21 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_41_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_203 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_23_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_92 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_70 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_47_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_38_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_429 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_204 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_590 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_82 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_71 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_60 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_93 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_63_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_47_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_419 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_56_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_3 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XTAP_205 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_591 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_94 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_83 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_72 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_61 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_50 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_409 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_30_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_206 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_592 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_95 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_84 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_73 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_62 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_40 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_51 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_43_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_207 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_593 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_33_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_390 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_96 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_85 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_74 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_63 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_41 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_52 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XANTENNA_output6_A x12/Y GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_18_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xx10 x9/B x2/A GND GND VDD VDD x12/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_208 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_43_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_41_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_17_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_561 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_594 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_391 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_20 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_31 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_42 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_97 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_86 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_75 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_361 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xx11 x4/X x6/B GND GND VDD VDD x12/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_62_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_209 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_25_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_584 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_595 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_392 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_98 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_87 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_76 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_65 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_21 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_32 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_43 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_54 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_55_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
Xx12 x12/A x12/B GND GND VDD VDD x12/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_38_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_18_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_20_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_596 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_393 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_88 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_77 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_66 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_22 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_33 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_44 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_55 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_33_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_190 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_55_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_18_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_24_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_597 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_520 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_350 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_394 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_89 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_78 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_67 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_23 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_34 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_45 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_56 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_59_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_41_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_180 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_191 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_59_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_44_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_16_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_543 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_598 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_384 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_395 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_24 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_35 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_46 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_79 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_68 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_57 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_181 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XANTENNA_x6_A x6/A GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_49_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_57_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_52_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_566 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_522 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_588 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_21 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_396 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_330 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_58 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_36 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_47 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_182 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_64_41 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_589 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_523 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_23 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_60_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_397 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_320 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_26 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_37 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_48 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_32_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_150 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_172 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_46_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_28_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_50_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_40_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_579 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_524 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_9 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_53_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_310 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_27 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_38 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_49 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_44_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_173 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_140 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_48_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_393 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_525 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_569 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_366 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_300 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_28 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XPHY_39 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_50_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_174 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_130 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_15_361 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_548 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_559 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_21_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_39_217 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_62_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_317 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_389 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_301 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_29 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xoutput4 x3/Y GND GND VDD VDD g0 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_109 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_186 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_13_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_51_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_549 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_321 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_42_26 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_38_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_41_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XTAP_379 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_44_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xoutput5 x9/Y GND GND VDD VDD g1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_132 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_49_335 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_64_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_64_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_265 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_385 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_539 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_12_333 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_303 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_44_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 GND GND VDD VDD sky130_ef_sc_hd__decap_12
Xoutput6 x12/Y GND GND VDD VDD rc sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 GND GND VDD VDD sky130_ef_sc_hd__decap_12
XTAP_166 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

