VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO encoder_proj
  CLASS BLOCK ;
  FOREIGN encoder_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END io_in[37]
  PIN io_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_in[38]
  PIN io_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_in[39]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END io_in[3]
  PIN io_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_in[40]
  PIN io_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END io_in[41]
  PIN io_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_in[42]
  PIN io_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_in[43]
  PIN io_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_in[44]
  PIN io_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_in[45]
  PIN io_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_in[46]
  PIN io_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END io_in[47]
  PIN io_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_in[48]
  PIN io_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END io_in[49]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END io_in[4]
  PIN io_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_in[50]
  PIN io_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END io_in[51]
  PIN io_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END io_in[52]
  PIN io_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_in[53]
  PIN io_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END io_in[54]
  PIN io_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_in[55]
  PIN io_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_in[56]
  PIN io_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END io_in[57]
  PIN io_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_in[58]
  PIN io_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_in[59]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_in[5]
  PIN io_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_in[60]
  PIN io_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[61]
  PIN io_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END io_in[62]
  PIN io_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END io_in[63]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 200.000 14.240 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 42.200 200.000 42.800 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.760 200.000 71.360 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 200.000 128.480 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 156.440 200.000 157.040 ;
    END
  END io_out[5]
  PIN valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.000 200.000 185.600 ;
    END
  END valid
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 4.690 10.695 192.650 187.865 ;
      LAYER met3 ;
        RECT 3.990 186.000 196.000 187.845 ;
        RECT 4.400 184.600 195.600 186.000 ;
        RECT 3.990 183.280 196.000 184.600 ;
        RECT 4.400 181.880 196.000 183.280 ;
        RECT 3.990 180.560 196.000 181.880 ;
        RECT 4.400 179.160 196.000 180.560 ;
        RECT 3.990 177.840 196.000 179.160 ;
        RECT 4.400 176.440 196.000 177.840 ;
        RECT 3.990 175.120 196.000 176.440 ;
        RECT 4.400 173.720 196.000 175.120 ;
        RECT 3.990 172.400 196.000 173.720 ;
        RECT 4.400 171.000 196.000 172.400 ;
        RECT 3.990 169.680 196.000 171.000 ;
        RECT 4.400 168.280 196.000 169.680 ;
        RECT 3.990 166.960 196.000 168.280 ;
        RECT 4.400 165.560 196.000 166.960 ;
        RECT 3.990 164.240 196.000 165.560 ;
        RECT 4.400 162.840 196.000 164.240 ;
        RECT 3.990 161.520 196.000 162.840 ;
        RECT 4.400 160.120 196.000 161.520 ;
        RECT 3.990 158.800 196.000 160.120 ;
        RECT 4.400 157.440 196.000 158.800 ;
        RECT 4.400 157.400 195.600 157.440 ;
        RECT 3.990 156.080 195.600 157.400 ;
        RECT 4.400 156.040 195.600 156.080 ;
        RECT 4.400 154.680 196.000 156.040 ;
        RECT 3.990 153.360 196.000 154.680 ;
        RECT 4.400 151.960 196.000 153.360 ;
        RECT 3.990 150.640 196.000 151.960 ;
        RECT 4.400 149.240 196.000 150.640 ;
        RECT 3.990 147.920 196.000 149.240 ;
        RECT 4.400 146.520 196.000 147.920 ;
        RECT 3.990 145.200 196.000 146.520 ;
        RECT 4.400 143.800 196.000 145.200 ;
        RECT 3.990 142.480 196.000 143.800 ;
        RECT 4.400 141.080 196.000 142.480 ;
        RECT 3.990 139.760 196.000 141.080 ;
        RECT 4.400 138.360 196.000 139.760 ;
        RECT 3.990 137.040 196.000 138.360 ;
        RECT 4.400 135.640 196.000 137.040 ;
        RECT 3.990 134.320 196.000 135.640 ;
        RECT 4.400 132.920 196.000 134.320 ;
        RECT 3.990 131.600 196.000 132.920 ;
        RECT 4.400 130.200 196.000 131.600 ;
        RECT 3.990 128.880 196.000 130.200 ;
        RECT 4.400 127.480 195.600 128.880 ;
        RECT 3.990 126.160 196.000 127.480 ;
        RECT 4.400 124.760 196.000 126.160 ;
        RECT 3.990 123.440 196.000 124.760 ;
        RECT 4.400 122.040 196.000 123.440 ;
        RECT 3.990 120.720 196.000 122.040 ;
        RECT 4.400 119.320 196.000 120.720 ;
        RECT 3.990 118.000 196.000 119.320 ;
        RECT 4.400 116.600 196.000 118.000 ;
        RECT 3.990 115.280 196.000 116.600 ;
        RECT 4.400 113.880 196.000 115.280 ;
        RECT 3.990 112.560 196.000 113.880 ;
        RECT 4.400 111.160 196.000 112.560 ;
        RECT 3.990 109.840 196.000 111.160 ;
        RECT 4.400 108.440 196.000 109.840 ;
        RECT 3.990 107.120 196.000 108.440 ;
        RECT 4.400 105.720 196.000 107.120 ;
        RECT 3.990 104.400 196.000 105.720 ;
        RECT 4.400 103.000 196.000 104.400 ;
        RECT 3.990 101.680 196.000 103.000 ;
        RECT 4.400 100.320 196.000 101.680 ;
        RECT 4.400 100.280 195.600 100.320 ;
        RECT 3.990 98.960 195.600 100.280 ;
        RECT 4.400 98.920 195.600 98.960 ;
        RECT 4.400 97.560 196.000 98.920 ;
        RECT 3.990 96.240 196.000 97.560 ;
        RECT 4.400 94.840 196.000 96.240 ;
        RECT 3.990 93.520 196.000 94.840 ;
        RECT 4.400 92.120 196.000 93.520 ;
        RECT 3.990 90.800 196.000 92.120 ;
        RECT 4.400 89.400 196.000 90.800 ;
        RECT 3.990 88.080 196.000 89.400 ;
        RECT 4.400 86.680 196.000 88.080 ;
        RECT 3.990 85.360 196.000 86.680 ;
        RECT 4.400 83.960 196.000 85.360 ;
        RECT 3.990 82.640 196.000 83.960 ;
        RECT 4.400 81.240 196.000 82.640 ;
        RECT 3.990 79.920 196.000 81.240 ;
        RECT 4.400 78.520 196.000 79.920 ;
        RECT 3.990 77.200 196.000 78.520 ;
        RECT 4.400 75.800 196.000 77.200 ;
        RECT 3.990 74.480 196.000 75.800 ;
        RECT 4.400 73.080 196.000 74.480 ;
        RECT 3.990 71.760 196.000 73.080 ;
        RECT 4.400 70.360 195.600 71.760 ;
        RECT 3.990 69.040 196.000 70.360 ;
        RECT 4.400 67.640 196.000 69.040 ;
        RECT 3.990 66.320 196.000 67.640 ;
        RECT 4.400 64.920 196.000 66.320 ;
        RECT 3.990 63.600 196.000 64.920 ;
        RECT 4.400 62.200 196.000 63.600 ;
        RECT 3.990 60.880 196.000 62.200 ;
        RECT 4.400 59.480 196.000 60.880 ;
        RECT 3.990 58.160 196.000 59.480 ;
        RECT 4.400 56.760 196.000 58.160 ;
        RECT 3.990 55.440 196.000 56.760 ;
        RECT 4.400 54.040 196.000 55.440 ;
        RECT 3.990 52.720 196.000 54.040 ;
        RECT 4.400 51.320 196.000 52.720 ;
        RECT 3.990 50.000 196.000 51.320 ;
        RECT 4.400 48.600 196.000 50.000 ;
        RECT 3.990 47.280 196.000 48.600 ;
        RECT 4.400 45.880 196.000 47.280 ;
        RECT 3.990 44.560 196.000 45.880 ;
        RECT 4.400 43.200 196.000 44.560 ;
        RECT 4.400 43.160 195.600 43.200 ;
        RECT 3.990 41.840 195.600 43.160 ;
        RECT 4.400 41.800 195.600 41.840 ;
        RECT 4.400 40.440 196.000 41.800 ;
        RECT 3.990 39.120 196.000 40.440 ;
        RECT 4.400 37.720 196.000 39.120 ;
        RECT 3.990 36.400 196.000 37.720 ;
        RECT 4.400 35.000 196.000 36.400 ;
        RECT 3.990 33.680 196.000 35.000 ;
        RECT 4.400 32.280 196.000 33.680 ;
        RECT 3.990 30.960 196.000 32.280 ;
        RECT 4.400 29.560 196.000 30.960 ;
        RECT 3.990 28.240 196.000 29.560 ;
        RECT 4.400 26.840 196.000 28.240 ;
        RECT 3.990 25.520 196.000 26.840 ;
        RECT 4.400 24.120 196.000 25.520 ;
        RECT 3.990 22.800 196.000 24.120 ;
        RECT 4.400 21.400 196.000 22.800 ;
        RECT 3.990 20.080 196.000 21.400 ;
        RECT 4.400 18.680 196.000 20.080 ;
        RECT 3.990 17.360 196.000 18.680 ;
        RECT 4.400 15.960 196.000 17.360 ;
        RECT 3.990 14.640 196.000 15.960 ;
        RECT 4.400 13.240 195.600 14.640 ;
        RECT 3.990 10.715 196.000 13.240 ;
  END
END encoder_proj
END LIBRARY

