magic
tech sky130A
magscale 1 2
timestamp 1727964749
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 38824 37584
<< obsm2 >>
rect 938 2139 38530 37573
<< metal3 >>
rect 39200 36184 40000 36304
rect 0 33192 800 33312
rect 39200 29656 40000 29776
rect 39200 23128 40000 23248
rect 0 19864 800 19984
rect 39200 16600 40000 16720
rect 39200 10072 40000 10192
rect 0 6536 800 6656
rect 39200 3544 40000 3664
<< obsm3 >>
rect 800 36384 39200 37569
rect 800 36104 39120 36384
rect 800 33392 39200 36104
rect 880 33112 39200 33392
rect 800 29856 39200 33112
rect 800 29576 39120 29856
rect 800 23328 39200 29576
rect 800 23048 39120 23328
rect 800 20064 39200 23048
rect 880 19784 39200 20064
rect 800 16800 39200 19784
rect 800 16520 39120 16800
rect 800 10272 39200 16520
rect 800 9992 39120 10272
rect 800 6736 39200 9992
rect 880 6456 39200 6736
rect 800 3744 39200 6456
rect 800 3464 39120 3744
rect 800 2143 39200 3464
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 0 6536 800 6656 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 39200 23128 40000 23248 6 io_oeb[0]
port 4 nsew signal output
rlabel metal3 s 39200 29656 40000 29776 6 io_oeb[1]
port 5 nsew signal output
rlabel metal3 s 39200 36184 40000 36304 6 io_oeb[2]
port 6 nsew signal output
rlabel metal3 s 39200 3544 40000 3664 6 io_out[0]
port 7 nsew signal output
rlabel metal3 s 39200 10072 40000 10192 6 io_out[1]
port 8 nsew signal output
rlabel metal3 s 39200 16600 40000 16720 6 io_out[2]
port 9 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 487904
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/arbiter_proj/runs/24_10_03_16_11/results/signoff/arbiter_proj.magic.gds
string GDS_START 74806
<< end >>

