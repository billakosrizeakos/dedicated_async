magic
tech sky130A
magscale 1 2
timestamp 1726499675
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 2128 558808 349840
<< obsm2 >>
rect 938 2139 558514 349829
<< metal3 >>
rect 0 338920 800 339040
rect 559200 338920 560000 339040
rect 0 317160 800 317280
rect 559200 317160 560000 317280
rect 0 295400 800 295520
rect 559200 295400 560000 295520
rect 0 273640 800 273760
rect 559200 273640 560000 273760
rect 0 251880 800 252000
rect 559200 251880 560000 252000
rect 0 230120 800 230240
rect 559200 230120 560000 230240
rect 0 208360 800 208480
rect 559200 208360 560000 208480
rect 0 186600 800 186720
rect 559200 186600 560000 186720
rect 0 164840 800 164960
rect 559200 164840 560000 164960
rect 0 143080 800 143200
rect 559200 143080 560000 143200
rect 0 121320 800 121440
rect 559200 121320 560000 121440
rect 0 99560 800 99680
rect 559200 99560 560000 99680
rect 0 77800 800 77920
rect 559200 77800 560000 77920
rect 0 56040 800 56160
rect 559200 56040 560000 56160
rect 0 34280 800 34400
rect 559200 34280 560000 34400
rect 0 12520 800 12640
rect 559200 12520 560000 12640
<< obsm3 >>
rect 798 339120 559200 349825
rect 880 338840 559120 339120
rect 798 317360 559200 338840
rect 880 317080 559120 317360
rect 798 295600 559200 317080
rect 880 295320 559120 295600
rect 798 273840 559200 295320
rect 880 273560 559120 273840
rect 798 252080 559200 273560
rect 880 251800 559120 252080
rect 798 230320 559200 251800
rect 880 230040 559120 230320
rect 798 208560 559200 230040
rect 880 208280 559120 208560
rect 798 186800 559200 208280
rect 880 186520 559120 186800
rect 798 165040 559200 186520
rect 880 164760 559120 165040
rect 798 143280 559200 164760
rect 880 143000 559120 143280
rect 798 121520 559200 143000
rect 880 121240 559120 121520
rect 798 99760 559200 121240
rect 880 99480 559120 99760
rect 798 78000 559200 99480
rect 880 77720 559120 78000
rect 798 56240 559200 77720
rect 880 55960 559120 56240
rect 798 34480 559200 55960
rect 880 34200 559120 34480
rect 798 12720 559200 34200
rect 880 12440 559120 12720
rect 798 2143 559200 12440
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal3 s 0 12520 800 12640 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 230120 800 230240 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 251880 800 252000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 273640 800 273760 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 295400 800 295520 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 317160 800 317280 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 338920 800 339040 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 186600 800 186720 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 208360 800 208480 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 559200 12520 560000 12640 6 io_out[0]
port 17 nsew signal output
rlabel metal3 s 559200 230120 560000 230240 6 io_out[10]
port 18 nsew signal output
rlabel metal3 s 559200 251880 560000 252000 6 io_out[11]
port 19 nsew signal output
rlabel metal3 s 559200 273640 560000 273760 6 io_out[12]
port 20 nsew signal output
rlabel metal3 s 559200 295400 560000 295520 6 io_out[13]
port 21 nsew signal output
rlabel metal3 s 559200 317160 560000 317280 6 io_out[14]
port 22 nsew signal output
rlabel metal3 s 559200 338920 560000 339040 6 io_out[15]
port 23 nsew signal output
rlabel metal3 s 559200 34280 560000 34400 6 io_out[1]
port 24 nsew signal output
rlabel metal3 s 559200 56040 560000 56160 6 io_out[2]
port 25 nsew signal output
rlabel metal3 s 559200 77800 560000 77920 6 io_out[3]
port 26 nsew signal output
rlabel metal3 s 559200 99560 560000 99680 6 io_out[4]
port 27 nsew signal output
rlabel metal3 s 559200 121320 560000 121440 6 io_out[5]
port 28 nsew signal output
rlabel metal3 s 559200 143080 560000 143200 6 io_out[6]
port 29 nsew signal output
rlabel metal3 s 559200 164840 560000 164960 6 io_out[7]
port 30 nsew signal output
rlabel metal3 s 559200 186600 560000 186720 6 io_out[8]
port 31 nsew signal output
rlabel metal3 s 559200 208360 560000 208480 6 io_out[9]
port 32 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 51676692
string GDS_FILE /home/vasilis/Internship/dedicated_async/openlane/user_proj/runs/24_09_16_17_04/results/signoff/user_proj.magic.gds
string GDS_START 180298
<< end >>

