VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO arbiter_proj
  CLASS BLOCK ;
  FOREIGN arbiter_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_in[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 115.640 200.000 116.240 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 200.000 148.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.920 200.000 181.520 ;
    END
  END io_oeb[2]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.720 200.000 18.320 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 50.360 200.000 50.960 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 83.000 200.000 83.600 ;
    END
  END io_out[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 4.690 10.695 192.650 187.865 ;
      LAYER met3 ;
        RECT 4.000 181.920 196.000 187.845 ;
        RECT 4.000 180.520 195.600 181.920 ;
        RECT 4.000 166.960 196.000 180.520 ;
        RECT 4.400 165.560 196.000 166.960 ;
        RECT 4.000 149.280 196.000 165.560 ;
        RECT 4.000 147.880 195.600 149.280 ;
        RECT 4.000 116.640 196.000 147.880 ;
        RECT 4.000 115.240 195.600 116.640 ;
        RECT 4.000 100.320 196.000 115.240 ;
        RECT 4.400 98.920 196.000 100.320 ;
        RECT 4.000 84.000 196.000 98.920 ;
        RECT 4.000 82.600 195.600 84.000 ;
        RECT 4.000 51.360 196.000 82.600 ;
        RECT 4.000 49.960 195.600 51.360 ;
        RECT 4.000 33.680 196.000 49.960 ;
        RECT 4.400 32.280 196.000 33.680 ;
        RECT 4.000 18.720 196.000 32.280 ;
        RECT 4.000 17.320 195.600 18.720 ;
        RECT 4.000 10.715 196.000 17.320 ;
  END
END arbiter_proj
END LIBRARY

